** Profile: "SCHEMATIC1-test1"  [ E:\LabADE\pg1-SCHEMATIC1-test1.sim ] 

** Creating circuit file "pg1-SCHEMATIC1-test1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10m 0 0.01m 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pg1-SCHEMATIC1.net" 


.END
