** Profile: "SCHEMATIC1-test2"  [ E:\LabADE\pg2-SCHEMATIC1-test2.sim ] 

** Creating circuit file "pg2-SCHEMATIC1-test2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 4m 0 0.01m SKIPBP 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pg2-SCHEMATIC1.net" 


.END
