** Profile: "SCHEMATIC1-test3"  [ E:\LabADE\pg3-SCHEMATIC1-test3.sim ] 

** Creating circuit file "pg3-SCHEMATIC1-test3.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100m 0 0.01m 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pg3-SCHEMATIC1.net" 


.END
